library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- display.vhd
-- This entity implements the feature described in the video
-- https://www.youtube.com/watch?v=dLh1n2dErzE

-- The display on the Basys2 is common anode, so each segment 
-- is "active low", i.e. lighs up, when a zero is written to the corresponding
-- bit in seg_ca_o and/or seg_dp_o.
-- Likewise, the four anode signals are active low too.

entity display is

    generic (
                SIMULATION : boolean := false
            );
    port (
             -- Clock input from crystal (for delay)
             clk_i       : in  std_logic;

             -- Decimal value to convert
             value_i     : in  std_logic_vector (7 downto 0);
             two_comp_i  : in  std_logic;

             -- Output segment display
             seg_ca_o    : out std_logic_vector (6 downto 0);
             seg_dp_o    : out std_logic;
             seg_an_o    : out std_logic_vector (3 downto 0));

end display;

architecture Structural of display is
    function get_counter_size (simulation : boolean) return integer
    is
    begin
        if simulation then
            return 2;
        else
            return 15; -- 40 ns * 2^15 = 1.3 ms 
        end if;
            
    end function;

    constant COUNTER_SIZE : integer := get_counter_size(SIMULATION);

    signal segment : std_logic_vector(1 downto 0) := (others => '0');
    signal counter : std_logic_vector(COUNTER_SIZE-1 downto 0) :=
    (others => '0');

    constant DIG_0 : std_logic_vector (7 downto 0) := "11000000";
    constant DIG_1 : std_logic_vector (7 downto 0) := "11111001";
    constant DIG_2 : std_logic_vector (7 downto 0) := "10100100";
    constant DIG_3 : std_logic_vector (7 downto 0) := "10110000";
    constant DIG_4 : std_logic_vector (7 downto 0) := "10011001";
    constant DIG_5 : std_logic_vector (7 downto 0) := "10010010";
    constant DIG_6 : std_logic_vector (7 downto 0) := "10000010";
    constant DIG_7 : std_logic_vector (7 downto 0) := "11111000";
    constant DIG_8 : std_logic_vector (7 downto 0) := "10000000";
    constant DIG_9 : std_logic_vector (7 downto 0) := "10010000"; 
    constant BLANK : std_logic_vector (7 downto 0) := "11111111"; 
    constant NEGAT : std_logic_vector (7 downto 0) := "10111111"; 

    -- This holds the contents of the EEPROM with 11 address lines
    -- and 8 data lines.
    -- The data is generated by the short ruby script display.rb.
    type eeprom_type is array (0 to (2**11)-1) of std_logic_vector(7 downto 0);
    constant data : eeprom_type := (
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_3, DIG_3,
        DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3,
        DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4,
        DIG_4, DIG_4, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5,
        DIG_5, DIG_5, DIG_5, DIG_5, DIG_6, DIG_6, DIG_6, DIG_6,
        DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_7, DIG_7,
        DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7,
        DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8,
        DIG_8, DIG_8, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9,
        DIG_9, DIG_9, DIG_9, DIG_9, DIG_0, DIG_0, DIG_0, DIG_0,
        DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3,
        DIG_3, DIG_3, DIG_3, DIG_3, DIG_4, DIG_4, DIG_4, DIG_4,
        DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_5, DIG_5,
        DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5,
        DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_6,
        DIG_6, DIG_6, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7,
        DIG_7, DIG_7, DIG_7, DIG_7, DIG_8, DIG_8, DIG_8, DIG_8,
        DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_9, DIG_9,
        DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9,
        DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_0,
        DIG_0, DIG_0, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_3, DIG_3,
        DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3,
        DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4,
        DIG_4, DIG_4, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5,
        DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1, DIG_2, DIG_3,
        DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9, DIG_0, DIG_1,
        DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7, DIG_8, DIG_9,
        DIG_0, DIG_1, DIG_2, DIG_3, DIG_4, DIG_5, DIG_6, DIG_7,
        DIG_8, DIG_7, DIG_6, DIG_5, DIG_4, DIG_3, DIG_2, DIG_1,
        DIG_0, DIG_9, DIG_8, DIG_7, DIG_6, DIG_5, DIG_4, DIG_3,
        DIG_2, DIG_1, DIG_0, DIG_9, DIG_8, DIG_7, DIG_6, DIG_5,
        DIG_4, DIG_3, DIG_2, DIG_1, DIG_0, DIG_9, DIG_8, DIG_7,
        DIG_6, DIG_5, DIG_4, DIG_3, DIG_2, DIG_1, DIG_0, DIG_9,
        DIG_8, DIG_7, DIG_6, DIG_5, DIG_4, DIG_3, DIG_2, DIG_1,
        DIG_0, DIG_9, DIG_8, DIG_7, DIG_6, DIG_5, DIG_4, DIG_3,
        DIG_2, DIG_1, DIG_0, DIG_9, DIG_8, DIG_7, DIG_6, DIG_5,
        DIG_4, DIG_3, DIG_2, DIG_1, DIG_0, DIG_9, DIG_8, DIG_7,
        DIG_6, DIG_5, DIG_4, DIG_3, DIG_2, DIG_1, DIG_0, DIG_9,
        DIG_8, DIG_7, DIG_6, DIG_5, DIG_4, DIG_3, DIG_2, DIG_1,
        DIG_0, DIG_9, DIG_8, DIG_7, DIG_6, DIG_5, DIG_4, DIG_3,
        DIG_2, DIG_1, DIG_0, DIG_9, DIG_8, DIG_7, DIG_6, DIG_5,
        DIG_4, DIG_3, DIG_2, DIG_1, DIG_0, DIG_9, DIG_8, DIG_7,
        DIG_6, DIG_5, DIG_4, DIG_3, DIG_2, DIG_1, DIG_0, DIG_9,
        DIG_8, DIG_7, DIG_6, DIG_5, DIG_4, DIG_3, DIG_2, DIG_1,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_3, DIG_3,
        DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3,
        DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4,
        DIG_4, DIG_4, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5,
        DIG_5, DIG_5, DIG_5, DIG_5, DIG_6, DIG_6, DIG_6, DIG_6,
        DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_7, DIG_7,
        DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7,
        DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8,
        DIG_8, DIG_8, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9,
        DIG_9, DIG_9, DIG_9, DIG_9, DIG_0, DIG_0, DIG_0, DIG_0,
        DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_0, DIG_0, DIG_0, DIG_0, DIG_0,
        DIG_0, DIG_0, DIG_0, DIG_0, DIG_0, DIG_9, DIG_9, DIG_9,
        DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_9, DIG_8,
        DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8, DIG_8,
        DIG_8, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7, DIG_7,
        DIG_7, DIG_7, DIG_7, DIG_6, DIG_6, DIG_6, DIG_6, DIG_6,
        DIG_6, DIG_6, DIG_6, DIG_6, DIG_6, DIG_5, DIG_5, DIG_5,
        DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_5, DIG_4,
        DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4, DIG_4,
        DIG_4, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3, DIG_3,
        DIG_3, DIG_3, DIG_3, DIG_2, DIG_2, DIG_2, DIG_2, DIG_2,
        DIG_2, DIG_2, DIG_2, DIG_2, DIG_2, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, DIG_1,
        DIG_1, DIG_1, DIG_1, DIG_1, DIG_1, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK, BLANK,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT, NEGAT,
        others => BLANK);

    signal address    : std_logic_vector(10 downto 0);
    signal data_value : std_logic_vector (7 downto 0);

begin

    process (clk_i)
    begin
        if rising_edge(clk_i) then
            if counter = 0 then
                segment <= segment + 1;
            end if;
            counter <= counter + 1;
        end if;
    end process;

    address <= two_comp_i & segment & value_i;
    data_value <= data(conv_integer(address));

    seg_ca_o <= data_value(6 downto 0);
    seg_dp_o <= data_value(7);

    seg_an_o <= "1110" when segment = "00" else
                "1101" when segment = "01" else
                "1011" when segment = "10" else
                "0111" when segment = "11";

end Structural;

