library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package vga_bitmap_pkg is
    type vga_bitmap_t is array(0 to 255) of std_logic_vector(1 downto 0);

    constant vga_bitmap_0 : vga_bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","01","00","00","00","00","00","01","00","00","00","00",
        "00","00","00","00","00","00","01","00","00","00","01","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","01","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

    constant vga_bitmap_1 : vga_bitmap_t := (
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","01","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","01","00","00","00","00","00","00","00",
        "00","00","00","00","00","01","01","01","01","01","01","01","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00",
        "00","00","00","00","00","00","00","00","00","00","00","00","00","00","00","00");

end package vga_bitmap_pkg;

