library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- output.vhd
-- This entity implements the feature described in the video
-- https://www.youtube.com/watch?v=dLh1n2dErzE

-- The display on the Basys2 is common anode, so each segment 
-- is "active low", i.e. lighs up, when a zero is written to the corresponding
-- bit in seg_ca_o and/or seg_dp_o.
-- Likewise, the four anode signals are active low too.

entity output is

    generic (
                COUNTER_SIZE : integer := 15
            -- 40 ns * 2^15 = 1.3 ms
            );
    port (
             -- Clock input from crystal (for delay)
             clk_i       : in  std_logic;

             -- Decimal value to convert
             value_i     : in  std_logic_vector (7 downto 0);

             -- Output segment display
             seg_ca_o    : out std_logic_vector (6 downto 0);
             seg_dp_o    : out std_logic;
             seg_an_o    : out std_logic_vector (3 downto 0));

end output;

architecture Structural of output is
    signal segment : std_logic_vector(1 downto 0) := (others => '0');
    signal counter : std_logic_vector(COUNTER_SIZE-1 downto 0) :=
    (others => '0');

    -- This holds the contents of the EEPROM with 11 address lines
    -- and 8 data lines.
    -- The data is generated by the short ruby script output.rb.
    type eeprom_type is array (0 to (2**11)-1) of std_logic_vector(7 downto 0);
    constant data : eeprom_type := (

    "11000000", "11111001", "10100100", "10110000", "10011001", "10010010", "10000010", "11111000",
    "10000000", "10010000", "11000000", "11111001", "10100100", "10110000", "10011001", "10010010",
    "10000010", "11111000", "10000000", "10010000", "11000000", "11111001", "10100100", "10110000",
    "10011001", "10010010", "10000010", "11111000", "10000000", "10010000", "11000000", "11111001",
    "10100100", "10110000", "10011001", "10010010", "10000010", "11111000", "10000000", "10010000",
    "11000000", "11111001", "10100100", "10110000", "10011001", "10010010", "10000010", "11111000",
    "10000000", "10010000", "11000000", "11111001", "10100100", "10110000", "10011001", "10010010",
    "10000010", "11111000", "10000000", "10010000", "11000000", "11111001", "10100100", "10110000",
    "10011001", "10010010", "10000010", "11111000", "10000000", "10010000", "11000000", "11111001",
    "10100100", "10110000", "10011001", "10010010", "10000010", "11111000", "10000000", "10010000",
    "11000000", "11111001", "10100100", "10110000", "10011001", "10010010", "10000010", "11111000",
    "10000000", "10010000", "11000000", "11111001", "10100100", "10110000", "10011001", "10010010",
    "10000010", "11111000", "10000000", "10010000", "11000000", "11111001", "10100100", "10110000",
    "10011001", "10010010", "10000010", "11111000", "10000000", "10010000", "11000000", "11111001",
    "10100100", "10110000", "10011001", "10010010", "10000010", "11111000", "10000000", "10010000",
    "11000000", "11111001", "10100100", "10110000", "10011001", "10010010", "10000010", "11111000",
    "10000000", "10010000", "11000000", "11111001", "10100100", "10110000", "10011001", "10010010",
    "10000010", "11111000", "10000000", "10010000", "11000000", "11111001", "10100100", "10110000",
    "10011001", "10010010", "10000010", "11111000", "10000000", "10010000", "11000000", "11111001",
    "10100100", "10110000", "10011001", "10010010", "10000010", "11111000", "10000000", "10010000",
    "11000000", "11111001", "10100100", "10110000", "10011001", "10010010", "10000010", "11111000",
    "10000000", "10010000", "11000000", "11111001", "10100100", "10110000", "10011001", "10010010",
    "10000010", "11111000", "10000000", "10010000", "11000000", "11111001", "10100100", "10110000",
    "10011001", "10010010", "10000010", "11111000", "10000000", "10010000", "11000000", "11111001",
    "10100100", "10110000", "10011001", "10010010", "10000010", "11111000", "10000000", "10010000",
    "11000000", "11111001", "10100100", "10110000", "10011001", "10010010", "10000010", "11111000",
    "10000000", "10010000", "11000000", "11111001", "10100100", "10110000", "10011001", "10010010",
    "10000010", "11111000", "10000000", "10010000", "11000000", "11111001", "10100100", "10110000",
    "10011001", "10010010", "10000010", "11111000", "10000000", "10010000", "11000000", "11111001",
    "10100100", "10110000", "10011001", "10010010", "10000010", "11111000", "10000000", "10010000",
    "11000000", "11111001", "10100100", "10110000", "10011001", "10010010", "10000010", "11111000",
    "10000000", "10010000", "11000000", "11111001", "10100100", "10110000", "10011001", "10010010",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10110000", "10110000",
    "10110000", "10110000", "10110000", "10110000", "10110000", "10110000", "10110000", "10110000",
    "10011001", "10011001", "10011001", "10011001", "10011001", "10011001", "10011001", "10011001",
    "10011001", "10011001", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010",
    "10010010", "10010010", "10010010", "10010010", "10000010", "10000010", "10000010", "10000010",
    "10000010", "10000010", "10000010", "10000010", "10000010", "10000010", "11111000", "11111000",
    "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000",
    "10000000", "10000000", "10000000", "10000000", "10000000", "10000000", "10000000", "10000000",
    "10000000", "10000000", "10010000", "10010000", "10010000", "10010000", "10010000", "10010000",
    "10010000", "10010000", "10010000", "10010000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10110000", "10110000", "10110000", "10110000", "10110000", "10110000",
    "10110000", "10110000", "10110000", "10110000", "10011001", "10011001", "10011001", "10011001",
    "10011001", "10011001", "10011001", "10011001", "10011001", "10011001", "10010010", "10010010",
    "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010",
    "10000010", "10000010", "10000010", "10000010", "10000010", "10000010", "10000010", "10000010",
    "10000010", "10000010", "11111000", "11111000", "11111000", "11111000", "11111000", "11111000",
    "11111000", "11111000", "11111000", "11111000", "10000000", "10000000", "10000000", "10000000",
    "10000000", "10000000", "10000000", "10000000", "10000000", "10000000", "10010000", "10010000",
    "10010000", "10010000", "10010000", "10010000", "10010000", "10010000", "10010000", "10010000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10110000", "10110000",
    "10110000", "10110000", "10110000", "10110000", "10110000", "10110000", "10110000", "10110000",
    "10011001", "10011001", "10011001", "10011001", "10011001", "10011001", "10011001", "10011001",
    "10011001", "10011001", "10010010", "10010010", "10010010", "10010010", "10010010", "10010010",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000", "11000000",
    "11000000", "11000000", "11000000", "11000000", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001", "11111001",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100", "10100100",
    others => "11111111");

    signal address    : std_logic_vector(10 downto 0);
    signal data_value : std_logic_vector (7 downto 0);

begin

    process (clk_i)
    begin
        if rising_edge(clk_i) then
            if counter = 0 then
                segment <= segment + 1;
            end if;
            counter <= counter + 1;
        end if;
    end process;

    address <= "0" & segment & value_i;
    data_value <= data(conv_integer(address));

    seg_ca_o <= data_value(6 downto 0);
    seg_dp_o <= data_value(7);

    seg_an_o <= "1110" when segment = "00" else
                "1101" when segment = "01" else
                "1011" when segment = "10" else
                "0111" when segment = "11";

end Structural;

