library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package vga_bitmap_pkg is
    type vga_bitmap_t is array(0 to 255) of std_logic;

    constant vga_bitmap_0 : vga_bitmap_t := (
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0',
        '0','0','0','0','0','0','1','0','0','0','1','0','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','1','0','0','0','0','0','1','0','0','0','0',
        '0','0','0','0','0','0','1','0','0','0','1','0','0','0','0','0',
        '0','0','0','0','0','0','0','1','1','1','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');

    constant vga_bitmap_1 : vga_bitmap_t := (
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','1','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','1','1','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
        '0','0','0','0','0','1','1','1','1','1','1','1','0','0','0','0',
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
        '0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');

end package vga_bitmap_pkg;

